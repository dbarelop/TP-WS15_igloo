LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

ENTITY AD7782_tb IS
	-- empty
END AD7782_tb;

ARCHITECTURE verhalten OF AD7782_tb IS


END verhalten;