LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY AD7782CTRL IS
-- now empty
END AD7782CTRL;


ARCHITECTURE behaviour OF AD7782CTRL IS

END behaviour;